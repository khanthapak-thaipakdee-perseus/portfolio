library verilog;
use verilog.vl_types.all;
entity compare_2_vlg_vec_tst is
end compare_2_vlg_vec_tst;
