library verilog;
use verilog.vl_types.all;
entity compare_4_vlg_vec_tst is
end compare_4_vlg_vec_tst;
